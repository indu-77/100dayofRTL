module mux(i,s,d);
input [7:0]i;
input [2:0]s;
output d;
reg d;
always @(s)
begin
case(s)
3'b000: d=i[0];
3'b001: d=i[1];
3'b010: d=i[2];
3'b011: d=i[3];
3'b100: d=i[4];
3'b101: d=i[5];
3'b110: d=i[6];
3'b111: d=i[7];
default d=1'bz;
endcase 
end
endmodule

module mux_tb;
wire d;
reg [7:0]i;
reg [2:0]s;
assign i=8'b11011100;
mux m1(i,s,d);
integer j;
initial
begin
for(j=0;j<8;j=j+1)
begin
#2{s}=j;
end
end
endmodule

